module multaddsub_add_sign_7_6(input logic a,b,
                                output logic c);
 
    assign c = a ^ b;
endmodule