module compile_test(input logic a,b,
                                output logic c);
 
    assign c = a ^ b;
endmodule